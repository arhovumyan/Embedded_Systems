`ifndef DEFINITIONS_VH
`define DEFINITIONS_VH

`define BIT_WIDTH 16
`define RESULT_WIDTH (2*`BIT_WIDTH)

`endif
