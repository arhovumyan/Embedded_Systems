`ifndef MM_DEFINITIONS_VH
`define MM_DEFINITIONS_VH

`define FACTOR_WIDTH_DEFAULT  16
`define PRODUCT_WIDTH_DEFAULT (`FACTOR_WIDTH_DEFAULT * 2 + 2)

`endif
