`timescale 1ns / 1ps

`default_nettype none
`include "mm_definitions.vh"

module mm_testbench;

  localparam integer NBITS  = `FACTOR_WIDTH_DEFAULT;
  localparam integer RESULT_WIDTH = `PRODUCT_WIDTH_DEFAULT;
  
  reg signed [NBITS-1:0] A_11, A_12, A_13, A_21, A_22, A_23, A_31, A_32, A_33, B_11, B_21, B_31;
  
  wire signed [RESULT_WIDTH-1:0] C_11, C_21, C_31;
    
  top_matrix_multiplication
  #(
        .NBITS(NBITS),
        .RESULT_WIDTH(RESULT_WIDTH)
  )
  controller
  (
      .A_11(A_11),
      .A_12(A_12),
      .A_13(A_13),
      .A_21(A_21),
      .A_22(A_22),
      .A_23(A_23),
      .A_31(A_31),
      .A_32(A_32),
      .A_33(A_33),
      .B_11(B_11),
      .B_21(B_21),
      .B_31(B_31),
      
      .C_11(C_11),
      .C_21(C_21),
      .C_31(C_31) 
  );
  
  initial begin
  A_11 = 0;
  A_12 = 0;
  A_13 = 0;
  A_21 = 0;
  A_22 = 0;
  A_23 = 0;
  A_31 = 0;
  A_32 = 0;
  A_33 = 0;
  B_11 = 0;
  B_21 = 0;
  B_31 = 0;
  
  #20
  A_11 = -12345;
A_12 =  2468;
A_13 = -31000;
A_21 =  15874;
A_22 = -8765;
A_23 =  9999;
A_31 = -32768;
A_32 =  32767;
A_33 =  5432;
B_11 = -11111;
B_21 =  22222;
B_31 = -13579;
  
  #20
A_11 =  30500;
A_12 = -25000;
A_13 =  1234;
A_21 = -16384;
A_22 =  3276;
A_23 =  999;
A_31 =  2048;
A_32 = -3072;
A_33 =  16383;
B_11 =  10000;
B_21 = -20000;
B_31 =  30000;

  
  #20
  A_11 = -7654;
A_12 =  4321;
A_13 =  28765;
A_21 = -12000;
A_22 =  876;
A_23 = -22222;
A_31 =  17000;
A_32 = -31415;
A_33 =  28000;
B_11 = -3276;
B_21 =  15000;
B_31 =  27000;

  #20
  A_11 =  1111;
A_12 = -2222;
A_13 =  3333;
A_21 = -4444;
A_22 =  5555;
A_23 = -6666;
A_31 =  7777;
A_32 = -8888;
A_33 =  9999;
B_11 = -1234;
B_21 =  24680;
B_31 = -1357;
  
  #20
  A_11 =  31000;
A_12 = -15000;
A_13 =  500;
A_21 = -25000;
A_22 =  16384;
A_23 = -8192;
A_31 =  27000;
A_32 = -32760;
A_33 =  12000;
B_11 =  32767;
B_21 = -32768;
B_31 =  12345;
  
  $finish;
  
  end
  
endmodule
